-- demo_soc.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity demo_soc is
	port (
		clk_clk            : in    std_logic                     := '0';             --    clk.clk
		memory_mem_a       : out   std_logic_vector(12 downto 0);                    -- memory.mem_a
		memory_mem_ba      : out   std_logic_vector(2 downto 0);                     --       .mem_ba
		memory_mem_ck      : out   std_logic;                                        --       .mem_ck
		memory_mem_ck_n    : out   std_logic;                                        --       .mem_ck_n
		memory_mem_cke     : out   std_logic;                                        --       .mem_cke
		memory_mem_cs_n    : out   std_logic;                                        --       .mem_cs_n
		memory_mem_ras_n   : out   std_logic;                                        --       .mem_ras_n
		memory_mem_cas_n   : out   std_logic;                                        --       .mem_cas_n
		memory_mem_we_n    : out   std_logic;                                        --       .mem_we_n
		memory_mem_reset_n : out   std_logic;                                        --       .mem_reset_n
		memory_mem_dq      : inout std_logic_vector(7 downto 0)  := (others => '0'); --       .mem_dq
		memory_mem_dqs     : inout std_logic                     := '0';             --       .mem_dqs
		memory_mem_dqs_n   : inout std_logic                     := '0';             --       .mem_dqs_n
		memory_mem_odt     : out   std_logic;                                        --       .mem_odt
		memory_mem_dm      : out   std_logic;                                        --       .mem_dm
		memory_oct_rzqin   : in    std_logic                     := '0';             --       .oct_rzqin
		reset_reset_n      : in    std_logic                     := '0'              --  reset.reset_n
	);
end entity demo_soc;

architecture rtl of demo_soc is
	component clk_gen_wrapper is
		port (
			rsi_rstn      : in  std_logic                     := 'X';             -- reset_n
			csi_clk       : in  std_logic                     := 'X';             -- clk
			trig_out      : out std_logic;                                        -- new_signal
			clk_out       : out std_logic;                                        -- clk
			avs_write     : in  std_logic                     := 'X';             -- write
			avs_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata  : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component clk_gen_wrapper;

	component dct_2d_ip_wrapper is
		port (
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_rstn        : in  std_logic                     := 'X';             -- reset_n
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dct_done        : out std_logic;                                        -- new_signal
			busy            : out std_logic;                                        -- new_signal
			start_dct       : in  std_logic                     := 'X';             -- new_signal
			new_output      : out std_logic;                                        -- new_signal
			new_output_data : out std_logic_vector(31 downto 0)                     -- new_signal
		);
	end component dct_2d_ip_wrapper;

	component delta_timer_wrapper is
		generic (
			REG_LAYER : boolean := false;
			CW        : integer := 7
		);
		port (
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_rstn        : in  std_logic                     := 'X';             -- reset_n
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			trig_in         : in  std_logic                     := 'X';             -- new_signal
			signal_from_DUV : in  std_logic                     := 'X';             -- new_signal
			trig_out        : out std_logic                                         -- new_signal
		);
	end component delta_timer_wrapper;

	component fifo_snk_wrapper is
		generic (
			DEPTH : integer := 8;
			DW    : integer := 32
		);
		port (
			csi_clk        : in  std_logic                     := 'X';             -- clk
			rsi_rstn       : in  std_logic                     := 'X';             -- reset_n
			avs_read       : in  std_logic                     := 'X';             -- read
			avs_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			avs_write      : in  std_logic                     := 'X';             -- write
			avs_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			trig_out       : out std_logic;                                        -- new_signal
			full_to_DUV    : out std_logic;                                        -- new_signal
			wr_from_DUV    : in  std_logic                     := 'X';             -- new_signal
			wdata_from_DUV : in  std_logic_vector(31 downto 0) := (others => 'X')  -- new_signal
		);
	end component fifo_snk_wrapper;

	component demo_soc_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a          : out   std_logic_vector(12 downto 0);                    -- mem_a
			mem_ba         : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck         : out   std_logic;                                        -- mem_ck
			mem_ck_n       : out   std_logic;                                        -- mem_ck_n
			mem_cke        : out   std_logic;                                        -- mem_cke
			mem_cs_n       : out   std_logic;                                        -- mem_cs_n
			mem_ras_n      : out   std_logic;                                        -- mem_ras_n
			mem_cas_n      : out   std_logic;                                        -- mem_cas_n
			mem_we_n       : out   std_logic;                                        -- mem_we_n
			mem_reset_n    : out   std_logic;                                        -- mem_reset_n
			mem_dq         : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs        : inout std_logic                     := 'X';             -- mem_dqs
			mem_dqs_n      : inout std_logic                     := 'X';             -- mem_dqs_n
			mem_odt        : out   std_logic;                                        -- mem_odt
			mem_dm         : out   std_logic;                                        -- mem_dm
			oct_rzqin      : in    std_logic                     := 'X';             -- oct_rzqin
			h2f_rst_n      : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID    : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR  : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN   : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE  : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK  : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT  : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID     : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA   : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB   : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST   : out   std_logic;                                        -- wlast
			h2f_lw_WVALID  : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY  : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID  : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY  : out   std_logic;                                        -- bready
			h2f_lw_ARID    : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR  : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN   : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE  : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK  : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT  : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST   : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID  : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY  : out   std_logic                                         -- rready
		);
	end component demo_soc_hps_0;

	component mode_selector_wrapper is
		port (
			csi_clk       : in  std_logic                     := 'X';             -- clk
			rsi_rstn      : in  std_logic                     := 'X';             -- reset_n
			avs_write     : in  std_logic                     := 'X';             -- write
			avs_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			mode_sel      : out std_logic                                         -- new_signal
		);
	end component mode_selector_wrapper;

	component re_det_wrapper is
		generic (
			REG_LAYER : boolean := false
		);
		port (
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_rstn        : in  std_logic                     := 'X';             -- reset_n
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			trig_out        : out std_logic;                                        -- new_signal
			signal_from_DUV : in  std_logic                     := 'X'              -- new_signal
		);
	end component re_det_wrapper;

	component rstn_gen_wrapper is
		generic (
			REG_LAYER : boolean := false
		);
		port (
			csi_clk         : in  std_logic                     := 'X';             -- clk
			rsi_rstn        : in  std_logic                     := 'X';             -- reset_n
			rso_rstn_to_DUV : out std_logic;                                        -- reset_n
			avs_write       : in  std_logic                     := 'X';             -- write
			avs_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			trig_out        : out std_logic                                         -- new_signal
		);
	end component rstn_gen_wrapper;

	component demo_soc_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			clk_gen_0_clk_out_clk                                               : in  std_logic                     := 'X';             -- clk
			clk_gen_0_reset_reset_bridge_in_reset_reset                         : in  std_logic                     := 'X';             -- reset
			delta_timer_0_reset_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			clk_gen_0_AVS_write                                                 : out std_logic;                                        -- write
			clk_gen_0_AVS_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			clk_gen_0_AVS_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			dct_2d_ip_0_avalon_slave_0_write                                    : out std_logic;                                        -- write
			dct_2d_ip_0_avalon_slave_0_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			delta_timer_0_AVS_write                                             : out std_logic;                                        -- write
			delta_timer_0_AVS_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			delta_timer_0_AVS_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_snk_0_avalon_slave_0_write                                     : out std_logic;                                        -- write
			fifo_snk_0_avalon_slave_0_read                                      : out std_logic;                                        -- read
			fifo_snk_0_avalon_slave_0_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_snk_0_avalon_slave_0_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			mode_selector_0_avalon_slave_0_write                                : out std_logic;                                        -- write
			mode_selector_0_avalon_slave_0_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mode_selector_0_avalon_slave_0_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			re_det_0_avalon_slave_0_write                                       : out std_logic;                                        -- write
			re_det_0_avalon_slave_0_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			re_det_0_avalon_slave_0_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			rstn_gen_0_AVS_write                                                : out std_logic;                                        -- write
			rstn_gen_0_AVS_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			rstn_gen_0_AVS_writedata                                            : out std_logic_vector(31 downto 0)                     -- writedata
		);
	end component demo_soc_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal clk_gen_0_clk_out_clk                                      : std_logic;                     -- clk_gen_0:clk_out -> [dct_2d_ip_0:csi_clk, delta_timer_0:csi_clk, fifo_snk_0:csi_clk, mm_interconnect_0:clk_gen_0_clk_out_clk, mode_selector_0:csi_clk, re_det_0:csi_clk, rst_controller_001:clk]
	signal dct_2d_ip_0_busy_new_signal                                : std_logic;                     -- dct_2d_ip_0:busy -> delta_timer_0:signal_from_DUV
	signal dct_2d_ip_0_new_output_new_signal                          : std_logic;                     -- dct_2d_ip_0:new_output -> fifo_snk_0:wr_from_DUV
	signal dct_2d_ip_0_dct_done_new_signal                            : std_logic;                     -- dct_2d_ip_0:dct_done -> re_det_0:signal_from_DUV
	signal mode_selector_0_mode_sel_new_signal                        : std_logic;                     -- mode_selector_0:mode_sel -> dct_2d_ip_0:start_dct
	signal dct_2d_ip_0_new_output_data_new_signal                     : std_logic_vector(31 downto 0); -- dct_2d_ip_0:new_output_data -> fifo_snk_0:wdata_from_DUV
	signal hps_0_h2f_lw_axi_master_awburst                            : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                              : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                              : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                             : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                             : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                              : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                            : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                             : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                             : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                             : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                             : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                              : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                            : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                            : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                               : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                             : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                             : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                             : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                            : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                            : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                            : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                             : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                             : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                              : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                              : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                               : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                             : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                             : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                            : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                             : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_delta_timer_0_avs_readdata               : std_logic_vector(31 downto 0); -- delta_timer_0:avs_readdata -> mm_interconnect_0:delta_timer_0_AVS_readdata
	signal mm_interconnect_0_delta_timer_0_avs_write                  : std_logic;                     -- mm_interconnect_0:delta_timer_0_AVS_write -> delta_timer_0:avs_write
	signal mm_interconnect_0_delta_timer_0_avs_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:delta_timer_0_AVS_writedata -> delta_timer_0:avs_writedata
	signal mm_interconnect_0_clk_gen_0_avs_readdata                   : std_logic_vector(31 downto 0); -- clk_gen_0:avs_readdata -> mm_interconnect_0:clk_gen_0_AVS_readdata
	signal mm_interconnect_0_clk_gen_0_avs_write                      : std_logic;                     -- mm_interconnect_0:clk_gen_0_AVS_write -> clk_gen_0:avs_write
	signal mm_interconnect_0_clk_gen_0_avs_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:clk_gen_0_AVS_writedata -> clk_gen_0:avs_writedata
	signal mm_interconnect_0_rstn_gen_0_avs_readdata                  : std_logic_vector(31 downto 0); -- rstn_gen_0:avs_readdata -> mm_interconnect_0:rstn_gen_0_AVS_readdata
	signal mm_interconnect_0_rstn_gen_0_avs_write                     : std_logic;                     -- mm_interconnect_0:rstn_gen_0_AVS_write -> rstn_gen_0:avs_write
	signal mm_interconnect_0_rstn_gen_0_avs_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:rstn_gen_0_AVS_writedata -> rstn_gen_0:avs_writedata
	signal mm_interconnect_0_re_det_0_avalon_slave_0_readdata         : std_logic_vector(31 downto 0); -- re_det_0:avs_readdata -> mm_interconnect_0:re_det_0_avalon_slave_0_readdata
	signal mm_interconnect_0_re_det_0_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:re_det_0_avalon_slave_0_write -> re_det_0:avs_write
	signal mm_interconnect_0_re_det_0_avalon_slave_0_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:re_det_0_avalon_slave_0_writedata -> re_det_0:avs_writedata
	signal mm_interconnect_0_fifo_snk_0_avalon_slave_0_readdata       : std_logic_vector(31 downto 0); -- fifo_snk_0:avs_readdata -> mm_interconnect_0:fifo_snk_0_avalon_slave_0_readdata
	signal mm_interconnect_0_fifo_snk_0_avalon_slave_0_read           : std_logic;                     -- mm_interconnect_0:fifo_snk_0_avalon_slave_0_read -> fifo_snk_0:avs_read
	signal mm_interconnect_0_fifo_snk_0_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:fifo_snk_0_avalon_slave_0_write -> fifo_snk_0:avs_write
	signal mm_interconnect_0_fifo_snk_0_avalon_slave_0_writedata      : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_snk_0_avalon_slave_0_writedata -> fifo_snk_0:avs_writedata
	signal mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_write         : std_logic;                     -- mm_interconnect_0:dct_2d_ip_0_avalon_slave_0_write -> dct_2d_ip_0:avs_write
	signal mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:dct_2d_ip_0_avalon_slave_0_writedata -> dct_2d_ip_0:avs_writedata
	signal mm_interconnect_0_mode_selector_0_avalon_slave_0_readdata  : std_logic_vector(31 downto 0); -- mode_selector_0:avs_readdata -> mm_interconnect_0:mode_selector_0_avalon_slave_0_readdata
	signal mm_interconnect_0_mode_selector_0_avalon_slave_0_write     : std_logic;                     -- mm_interconnect_0:mode_selector_0_avalon_slave_0_write -> mode_selector_0:avs_write
	signal mm_interconnect_0_mode_selector_0_avalon_slave_0_writedata : std_logic_vector(31 downto 0); -- mm_interconnect_0:mode_selector_0_avalon_slave_0_writedata -> mode_selector_0:avs_writedata
	signal rst_controller_reset_out_reset                             : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:clk_gen_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                         : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:delta_timer_0_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rstn_gen_0_reset_source_reset                              : std_logic;                     -- rstn_gen_0:rso_rstn_to_DUV -> rstn_gen_0_reset_source_reset:in
	signal rst_controller_002_reset_out_reset                         : std_logic;                     -- rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal hps_0_h2f_reset_reset                                      : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal reset_reset_n_ports_inv                                    : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [clk_gen_0:rsi_rstn, rstn_gen_0:rsi_rstn]
	signal rst_controller_001_reset_out_reset_ports_inv               : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [dct_2d_ip_0:rsi_rstn, delta_timer_0:rsi_rstn, fifo_snk_0:rsi_rstn, mode_selector_0:rsi_rstn, re_det_0:rsi_rstn]
	signal rstn_gen_0_reset_source_reset_ports_inv                    : std_logic;                     -- rstn_gen_0_reset_source_reset:inv -> rst_controller_001:reset_in0
	signal hps_0_h2f_reset_reset_ports_inv                            : std_logic;                     -- hps_0_h2f_reset_reset:inv -> rst_controller_002:reset_in0

begin

	clk_gen_0 : component clk_gen_wrapper
		port map (
			rsi_rstn      => rst_controller_reset_out_reset_ports_inv,  --    reset.reset_n
			csi_clk       => clk_clk,                                   --    clock.clk
			trig_out      => open,                                      -- trig_out.new_signal
			clk_out       => clk_gen_0_clk_out_clk,                     --  clk_out.clk
			avs_write     => mm_interconnect_0_clk_gen_0_avs_write,     --      AVS.write
			avs_writedata => mm_interconnect_0_clk_gen_0_avs_writedata, --         .writedata
			avs_readdata  => mm_interconnect_0_clk_gen_0_avs_readdata   --         .readdata
		);

	dct_2d_ip_0 : component dct_2d_ip_wrapper
		port map (
			csi_clk         => clk_gen_0_clk_out_clk,                                  --           clock.clk
			rsi_rstn        => rst_controller_001_reset_out_reset_ports_inv,           --           reset.reset_n
			avs_write       => mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_write,     --  avalon_slave_0.write
			avs_writedata   => mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_writedata, --                .writedata
			dct_done        => dct_2d_ip_0_dct_done_new_signal,                        --        dct_done.new_signal
			busy            => dct_2d_ip_0_busy_new_signal,                            --            busy.new_signal
			start_dct       => mode_selector_0_mode_sel_new_signal,                    --       start_dct.new_signal
			new_output      => dct_2d_ip_0_new_output_new_signal,                      --      new_output.new_signal
			new_output_data => dct_2d_ip_0_new_output_data_new_signal                  -- new_output_data.new_signal
		);

	delta_timer_0 : component delta_timer_wrapper
		generic map (
			REG_LAYER => false,
			CW        => 20
		)
		port map (
			csi_clk         => clk_gen_0_clk_out_clk,                         --           clock.clk
			rsi_rstn        => rst_controller_001_reset_out_reset_ports_inv,  --           reset.reset_n
			avs_write       => mm_interconnect_0_delta_timer_0_avs_write,     --             AVS.write
			avs_writedata   => mm_interconnect_0_delta_timer_0_avs_writedata, --                .writedata
			avs_readdata    => mm_interconnect_0_delta_timer_0_avs_readdata,  --                .readdata
			trig_in         => open,                                          --         trig_in.new_signal
			signal_from_DUV => dct_2d_ip_0_busy_new_signal,                   -- signal_from_DUV.new_signal
			trig_out        => open                                           --        trig_out.new_signal
		);

	fifo_snk_0 : component fifo_snk_wrapper
		generic map (
			DEPTH => 64,
			DW    => 32
		)
		port map (
			csi_clk        => clk_gen_0_clk_out_clk,                                 --          clock.clk
			rsi_rstn       => rst_controller_001_reset_out_reset_ports_inv,          --          reset.reset_n
			avs_read       => mm_interconnect_0_fifo_snk_0_avalon_slave_0_read,      -- avalon_slave_0.read
			avs_readdata   => mm_interconnect_0_fifo_snk_0_avalon_slave_0_readdata,  --               .readdata
			avs_write      => mm_interconnect_0_fifo_snk_0_avalon_slave_0_write,     --               .write
			avs_writedata  => mm_interconnect_0_fifo_snk_0_avalon_slave_0_writedata, --               .writedata
			trig_out       => open,                                                  --       trig_out.new_signal
			full_to_DUV    => open,                                                  --    full_to_DUV.new_signal
			wr_from_DUV    => dct_2d_ip_0_new_output_new_signal,                     --    wr_from_DUV.new_signal
			wdata_from_DUV => dct_2d_ip_0_new_output_data_new_signal                 -- wdata_from_DUV.new_signal
		);

	hps_0 : component demo_soc_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a          => memory_mem_a,                    --            memory.mem_a
			mem_ba         => memory_mem_ba,                   --                  .mem_ba
			mem_ck         => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n       => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke        => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n       => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n      => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n      => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n       => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n    => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq         => memory_mem_dq,                   --                  .mem_dq
			mem_dqs        => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n      => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt        => memory_mem_odt,                  --                  .mem_odt
			mem_dm         => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin      => memory_oct_rzqin,                --                  .oct_rzqin
			h2f_rst_n      => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_lw_axi_clk => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID    => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR  => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN   => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE  => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK  => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT  => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID     => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA   => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB   => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST   => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID  => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY  => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID     => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP   => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID  => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY  => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID    => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR  => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN   => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE  => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK  => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT  => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID     => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA   => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP   => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST   => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID  => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY  => hps_0_h2f_lw_axi_master_rready   --                  .rready
		);

	mode_selector_0 : component mode_selector_wrapper
		port map (
			csi_clk       => clk_gen_0_clk_out_clk,                                      --          clock.clk
			rsi_rstn      => rst_controller_001_reset_out_reset_ports_inv,               --          reset.reset_n
			avs_write     => mm_interconnect_0_mode_selector_0_avalon_slave_0_write,     -- avalon_slave_0.write
			avs_writedata => mm_interconnect_0_mode_selector_0_avalon_slave_0_writedata, --               .writedata
			avs_readdata  => mm_interconnect_0_mode_selector_0_avalon_slave_0_readdata,  --               .readdata
			mode_sel      => mode_selector_0_mode_sel_new_signal                         --       mode_sel.new_signal
		);

	re_det_0 : component re_det_wrapper
		generic map (
			REG_LAYER => false
		)
		port map (
			csi_clk         => clk_gen_0_clk_out_clk,                               --           clock.clk
			rsi_rstn        => rst_controller_001_reset_out_reset_ports_inv,        --           reset.reset_n
			avs_write       => mm_interconnect_0_re_det_0_avalon_slave_0_write,     --  avalon_slave_0.write
			avs_writedata   => mm_interconnect_0_re_det_0_avalon_slave_0_writedata, --                .writedata
			avs_readdata    => mm_interconnect_0_re_det_0_avalon_slave_0_readdata,  --                .readdata
			trig_out        => open,                                                --        trig_out.new_signal
			signal_from_DUV => dct_2d_ip_0_dct_done_new_signal                      -- signal_from_DUV.new_signal
		);

	rstn_gen_0 : component rstn_gen_wrapper
		generic map (
			REG_LAYER => false
		)
		port map (
			csi_clk         => clk_clk,                                    --        clock.clk
			rsi_rstn        => rst_controller_reset_out_reset_ports_inv,   --        reset.reset_n
			rso_rstn_to_DUV => rstn_gen_0_reset_source_reset,              -- reset_source.reset_n
			avs_write       => mm_interconnect_0_rstn_gen_0_avs_write,     --          AVS.write
			avs_writedata   => mm_interconnect_0_rstn_gen_0_avs_writedata, --             .writedata
			avs_readdata    => mm_interconnect_0_rstn_gen_0_avs_readdata,  --             .readdata
			trig_out        => open                                        --     trig_out.new_signal
		);

	mm_interconnect_0 : component demo_soc_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                               --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                             --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                              --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                             --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                            --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                             --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                            --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                             --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                            --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                            --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                              --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                              --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                              --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                             --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                             --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                              --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                             --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                             --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                               --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                             --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                              --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                             --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                            --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                             --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                            --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                             --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                            --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                            --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                              --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                              --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                              --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                             --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                             --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                    --                                                     clk_0_clk.clk
			clk_gen_0_clk_out_clk                                               => clk_gen_0_clk_out_clk,                                      --                                             clk_gen_0_clk_out.clk
			clk_gen_0_reset_reset_bridge_in_reset_reset                         => rst_controller_reset_out_reset,                             --                         clk_gen_0_reset_reset_bridge_in_reset.reset
			delta_timer_0_reset_reset_bridge_in_reset_reset                     => rst_controller_001_reset_out_reset,                         --                     delta_timer_0_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                         -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			clk_gen_0_AVS_write                                                 => mm_interconnect_0_clk_gen_0_avs_write,                      --                                                 clk_gen_0_AVS.write
			clk_gen_0_AVS_readdata                                              => mm_interconnect_0_clk_gen_0_avs_readdata,                   --                                                              .readdata
			clk_gen_0_AVS_writedata                                             => mm_interconnect_0_clk_gen_0_avs_writedata,                  --                                                              .writedata
			dct_2d_ip_0_avalon_slave_0_write                                    => mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_write,         --                                    dct_2d_ip_0_avalon_slave_0.write
			dct_2d_ip_0_avalon_slave_0_writedata                                => mm_interconnect_0_dct_2d_ip_0_avalon_slave_0_writedata,     --                                                              .writedata
			delta_timer_0_AVS_write                                             => mm_interconnect_0_delta_timer_0_avs_write,                  --                                             delta_timer_0_AVS.write
			delta_timer_0_AVS_readdata                                          => mm_interconnect_0_delta_timer_0_avs_readdata,               --                                                              .readdata
			delta_timer_0_AVS_writedata                                         => mm_interconnect_0_delta_timer_0_avs_writedata,              --                                                              .writedata
			fifo_snk_0_avalon_slave_0_write                                     => mm_interconnect_0_fifo_snk_0_avalon_slave_0_write,          --                                     fifo_snk_0_avalon_slave_0.write
			fifo_snk_0_avalon_slave_0_read                                      => mm_interconnect_0_fifo_snk_0_avalon_slave_0_read,           --                                                              .read
			fifo_snk_0_avalon_slave_0_readdata                                  => mm_interconnect_0_fifo_snk_0_avalon_slave_0_readdata,       --                                                              .readdata
			fifo_snk_0_avalon_slave_0_writedata                                 => mm_interconnect_0_fifo_snk_0_avalon_slave_0_writedata,      --                                                              .writedata
			mode_selector_0_avalon_slave_0_write                                => mm_interconnect_0_mode_selector_0_avalon_slave_0_write,     --                                mode_selector_0_avalon_slave_0.write
			mode_selector_0_avalon_slave_0_readdata                             => mm_interconnect_0_mode_selector_0_avalon_slave_0_readdata,  --                                                              .readdata
			mode_selector_0_avalon_slave_0_writedata                            => mm_interconnect_0_mode_selector_0_avalon_slave_0_writedata, --                                                              .writedata
			re_det_0_avalon_slave_0_write                                       => mm_interconnect_0_re_det_0_avalon_slave_0_write,            --                                       re_det_0_avalon_slave_0.write
			re_det_0_avalon_slave_0_readdata                                    => mm_interconnect_0_re_det_0_avalon_slave_0_readdata,         --                                                              .readdata
			re_det_0_avalon_slave_0_writedata                                   => mm_interconnect_0_re_det_0_avalon_slave_0_writedata,        --                                                              .writedata
			rstn_gen_0_AVS_write                                                => mm_interconnect_0_rstn_gen_0_avs_write,                     --                                                rstn_gen_0_AVS.write
			rstn_gen_0_AVS_readdata                                             => mm_interconnect_0_rstn_gen_0_avs_readdata,                  --                                                              .readdata
			rstn_gen_0_AVS_writedata                                            => mm_interconnect_0_rstn_gen_0_avs_writedata                  --                                                              .writedata
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => rstn_gen_0_reset_source_reset_ports_inv, -- reset_in0.reset
			clk            => clk_gen_0_clk_out_clk,                   --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                    -- (terminated)
			reset_req_in0  => '0',                                     -- (terminated)
			reset_in1      => '0',                                     -- (terminated)
			reset_req_in1  => '0',                                     -- (terminated)
			reset_in2      => '0',                                     -- (terminated)
			reset_req_in2  => '0',                                     -- (terminated)
			reset_in3      => '0',                                     -- (terminated)
			reset_req_in3  => '0',                                     -- (terminated)
			reset_in4      => '0',                                     -- (terminated)
			reset_req_in4  => '0',                                     -- (terminated)
			reset_in5      => '0',                                     -- (terminated)
			reset_req_in5  => '0',                                     -- (terminated)
			reset_in6      => '0',                                     -- (terminated)
			reset_req_in6  => '0',                                     -- (terminated)
			reset_in7      => '0',                                     -- (terminated)
			reset_req_in7  => '0',                                     -- (terminated)
			reset_in8      => '0',                                     -- (terminated)
			reset_req_in8  => '0',                                     -- (terminated)
			reset_in9      => '0',                                     -- (terminated)
			reset_req_in9  => '0',                                     -- (terminated)
			reset_in10     => '0',                                     -- (terminated)
			reset_req_in10 => '0',                                     -- (terminated)
			reset_in11     => '0',                                     -- (terminated)
			reset_req_in11 => '0',                                     -- (terminated)
			reset_in12     => '0',                                     -- (terminated)
			reset_req_in12 => '0',                                     -- (terminated)
			reset_in13     => '0',                                     -- (terminated)
			reset_req_in13 => '0',                                     -- (terminated)
			reset_in14     => '0',                                     -- (terminated)
			reset_req_in14 => '0',                                     -- (terminated)
			reset_in15     => '0',                                     -- (terminated)
			reset_req_in15 => '0'                                      -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rstn_gen_0_reset_source_reset_ports_inv <= not rstn_gen_0_reset_source_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of demo_soc
